// Hello world from SV classes

class day22;

  function new();
    // Leave Empty
  endfunction

  function void hello();
    $display("MERL, 2022\n");
  endfunction

endclass